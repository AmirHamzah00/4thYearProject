module NeuralNetwork (input logic clk, reset,
                     output logic [3:0] n0_weights [3:0]);
							
			
							
endmodule 